的	白 勺
我	手 戈
你	亻 尔
是	日 𤴓
了	㇇ 亅
不	丆 卜
在	𠂇 亻 土
他	亻 也
們	亻 門
我們
好	女 子
有	𠂇 月
這	辶 言
會	亼 口 丨 丷 日
嗎	口 馬
什	亻 十
麼	麻 幺
什麼
說	言 兌
她	女 也
想	相 心
一	一
很	彳 艮
人	㇒
那	刀 二 阝
來	木 从
都	者 阝
個	亻 固
能	䏍 匕
去	土 厶
和	禾 口
做	亻 故
上	⺊ 一
沒	氵 ㇆ 又
沒有
看	龵 目
怎	乍 心
怎麼
現	王 見
現在
點	黑 占
呢	口 尼
太	大 丶
裡	衤 里
聽	耳 王 𢛳
誰	言 隹
多	夕
時	日 寺
候	亻 丨 ユ 矢 
時候
下	一 卜
謝	言 射
謝謝
先	⺧ 儿
生	龶 ㇒
先生
喜	士 口 丷 一 口
歡	雚 欠
喜歡
大	人 一
東	木 日
西	兀 囗
東西
小	亅 八
叫	口 丩
愛	爫 冖 心 夂
年	𠂉 㐄
請	言 青
回	囗
工	一 丄
作	亻 乍
工作
錢	金 戔
吃	口 乞
開	門 开
家	宀 豕
哪	口 那
朋	月
友	𠂇 又
朋友
媽	女 馬
媽媽
今	亽 ㇇
天	一 大
今天
幾	戈 幺 
爸	父 巴
爸爸
些	此 二
樣	木 羕
怎麼樣
對	丷 一 羊 寸
起	走 己
對不起
住	亻 主
三	一 二
高	亠 口 冋
興	臼 冂 一 口 一 八
高興
買	罒 貝
醫	殹 酉
醫生
兒	臼 儿
哪兒
字	宀 子
名	夕 口
名字
認	言 忍
識	言 音 戈
認識
坐	土 从
喝	口 曷
寫	宀 舄
月	冂 二
號	号 虎
狗	犭 句
歲	止 厂 戈 一 小 丿
見	目 儿
看見
打	扌 丁
電	雨 电
話	言 舌
打電話
喂	口 畏
子	了 一
兒子
漂	氵 票
亮	亠 口 冖 几
漂亮
分	八 刀
鐘	金 童
分鐘
再	一 冉
再見
本	木 一
明	日 月
明天
少	小 丿
多少
塊	土 鬼
女	㇛ 丆
女兒
姐	女 且
小姐
衣	亠 𧘇
服	月 𠬝
衣服
水	水
學	𦥯 子
校	木 交
學校
影	景 彡
電影
書	聿 日
四	囗 儿
五	一 力 一
院	阝 完
醫院
關	門 幺 關
系	㇒ 糸
沒關系
飛	升
機	木 幾
飛機
二	一
視	礻 見
電視
讀	言 賣
後	彳 幺 夂
面	丆 囬
後面
昨	日 乍
昨天
睡	目 垂
覺	𦥯 見
睡覺
六	亠 八
老	耂 匕
師	𠂤 帀
老師
星	日 生
期	其 月
星期
十	一 丨
貓	豸 苗
腦	月 巛 囗 丶 乂
電腦
熱	埶 灬
學生
午	干 ㇒
下午
習	羽 白
學習
冷	冫 令
客	宀 各
氣	气 米
不客氣
前	䒑 刖
前面
八	㇒
中	口 丨
國	囗 或
中國
七	乚 一
菜	艹 采
桌	⺊ 日 木
桌子
出	山
租	禾 且
車	二 丨 日
出租車
天氣
茶	艹 人 十 八
九	丿 ㇈
商	亠 丷 冏
店	广 占
商店
椅	木 奇
椅子
同	冂 一 口
同學
一點
蘋	艹 頻
果	田 木
蘋果
飯	飠 反
飯店
中午
上午
水果
杯	木 不
杯子
雨	帀 冫
下雨
米	木 丷
米飯
北	匕
京	亠 口 小
北京
漢	氵 艹 口 丨 人 二
語	言 吾
漢語
就	京 尤
要	覀 女
知	矢 口
道	辶 首
知道
吧	口 巴
到	至 刂
也	乚 ㇆ 丨
還	辶 睘
讓	言 襄
給	糹 合
過	辶 咼
得	彳 㝵
真	十 具
著	艹 者
可	丁 口
以	乚 丶 人
可以
別	口 丿 ㇆ 刂
走	土 龰
告	⺧ 口
訴	言 斥
告訴
因	囗 大
為	丿 丶 ㇆ 灬
因為
快	忄 夬
但	亻 旦
但是
已	己
經	糹 巠
已經
為什麼
覺得
它	宀 匕
從	彳 从 龰
找	扌 戈
最	曰 取
可能
次	冫 欠
孩	子 亥
孩子
所	戶 斤
所以
兩	一 巾 从
錯	金 昔
等	⺮ 寺
題	是 頁
問	門 口
問題
一起
始	女 台
開始
間	門 日
時間
事	十 口 丨 ⺺ 亅
情	忄 青
事情
一下
非	非
常	龸 吊
非常
希	乂 布
望	肓 王
希望
準	淮 十
備	亻 艹 厂 用
準備
比	匕
件	亻 牛
意	音 心
思	田 心
意思
第	⺮ 弓 丨 ㇒
第一
進	辶 隹
大家
新	亲 斤
您	你 心
穿	穴 牙
送	辶 关
玩	王 元
長
小時
完	宀 元
每	𠂉 母
公	八 厶
司	㇆ 一 口
公司
幫	封 帛
助	且 力
幫助
晚	日 免
晚上
說話
門
忙	忄 亡
賣	士 罒 貝
房	户 方
房間
路	⻊ 各
懂	忄 董
正	一 止
正在
笑	⺮ 夭
遠	辶 袁
妻	十 ⺺ 女
妻子
丈	十 乂
夫	人 二
丈夫
離	离 隹
往	彳 主
男	田 力
眼	目 艮
睛	目 青
眼睛
樂	白 幺 木 
快樂
雖	虽 隹
然	肰 灬
雖然
早	日 十
早上
藥	艹 樂
身	㇆ 丨 ㇒ 二 丿
體	骨 豊
身體
黑
咖	口 加
啡	口 非
咖啡
日	口 一
休	亻 木
息	自 心
休息
外	夕 卜
生日
哥	可
哥哥
票	覀 示
手	㇒ 扌
手機
洗	氵 先
跳	⻊ 兆
舞	𠂉 卌 一 舛
跳舞
弟	丷 弓 丿 丨
弟弟
妹	女 未
妹妹
紅	糹 工
慢	忄 曼
近	辶 斤
白	日 ㇒
姐姐
介	人 丿 丨
紹	糹 召
介紹
魚	⺈ 田 灬
累	田 糸
課	言 果
班	玨 丿 丶
上班
旁	亠 丷 冖 方
邊	辶 臱
旁邊
運	辶 軍
動	重 力
運動
去年
報	幸 𠬝
紙	糹 氏
報紙
顏	彥 頁
色	⺈ 巴
顏色
場	土 昜
機場
唱	口 昌
歌	哥 欠
唱歌
千	㇒ 十
好吃
考	耂 丂
試	言 式
考試
左	𠂇 工
左邊
姓	女 生
百	一 白
雪	雨 彐
貴	中 一 貝
病	疒 丙
生病
游	氵 斿
泳	氵 永
游泳
牛	牛
奶	女 乃
牛奶
右	𠂇 口
右邊
便	亻 更
宜	宀 且
便宜
共	龷 八
汽	氵 气
公共汽車
床	广 木
起床
籃	⺮ 監
球	王 求
打籃球
雞	奚 隹
蛋	疋 虫
雞蛋
踢	⻊ 易
足	口 龰
踢足球
零	雨 令
表	龶 𧘇
手表
旅	方 丿 一 氏
旅游
務	矛 务
員	口 貝
服務員
賓	宀 一 小 丿 貝
館	飠 官
賓館
教	孝 ⺙
室	宀 至
教室
跑	⻊ 包
步	止 小 丿
跑步
陰	阝 侌
條	亻 丨 条
面條
鉛	金 几 口
筆	⺮ 聿
鉛筆
火  人 ㇒
站	立 占
火車站
瓜
西瓜
羊
肉	仌 冂
羊肉
晴	日 青
啊	口 阿
把	扌 巴
如	女 口
如果
只	口 八
被	衤 皮
跟	⻊ 艮
自	目 丶
己
自己
用
像	亻 象
需	雨 而
需要
應	䧹 心
該	言 亥
應該
起來
才	𠂇 ㇒
又	㇇ ㇏
拿	合 手
更	一 日 丨 乂
帶	儿 廿 冖 巾
然後
一樣
當	⺌ 冖 口 田
當然
相	木 目
信	亻 言
相信
認為
明白
直	十 目 一
一直
地	土 也
方
地方
離開
定	宀 𤴓
一定
還是
發	癶 弓 殳
發現
而	丆 𦉫
且	月 一
而且
必	心 丿
須	彡 頁
必須
放	方 ⺙
為了
向	宀 口
位	亻 立
種	禾 重
后	⺁ 一 口
最后
其	甘 一 八
其他
記	言 几
記得
或	戓 一
者	耂 日
或者
過去
擔	扌 詹
心	㇃ 丶
擔心
以前
世	㇗ 廿
界	田 介
世界
重	千 里
重要
別人
機會
張	弓 長
接	扌 妾
賽	宀 二 一 八 貝
比賽
關系
馬	一 二 丨 ㇉ 灬
馬上
決	氵 夬
決定
於	方 仒
關於
難	口 夫 廿 隹
瞭	目 尞
解	角 刀 牛
瞭解
結	糹 吉
束	木 口
結束
清	氵 青
楚	林 疋
清楚
願	原 頁
願意
花	艹 化
照	昭 灬
片  丿 丄 ㇕
照片
迎	辶 卬
歡迎
總	糹 悤
總是
嘴	口 觜
參	厽 㐱
加	力 口
參加
辦	辡 力
法	氵 去
辦法
選	辶 巽
擇	扌 睪
選擇
壞	土 褱
算	⺮ 目 一 丿 丨
打算
特	牛 寺
特別
注	氵 主
注意
實	宀 貫
其實
小心
久	勹 ㇏
只有
講	言 冓
故	古 ⺙
故事
換	扌 奐
婚	女 昏
結婚
段	丨 ㇒ 二 一 殳
努	奴 力
力	㇆ 丿
努力
害  宀 丄 二 口
怕	忄 白
害怕
剛	岡 刂
剛才
節	⺮ 即
目	口 二
節目
輛	車 兩
萬	艹 禺
解決
辦公室
奇	大 可
怪	忄 圣
奇怪
同意
戲	䖒 戈
游戲
幫忙
國家
最近
聲	殸 耳
音	立 日
聲音
可愛
成	万 戈
完成
半	二 丨 丷
求	𠂇 丶 氺
要求
除	阝 余
除了
容	宀 谷
易	日 勿
容易
臉	月 僉
簡	⺮ 間
單	吅 田 十
簡單
檢	木 僉
查	木 旦
檢查
音樂
越	走 戉
顧	雇 頁
照顧
聰	耳 悤
聰明
甜	舌 甘
突	穴 犬
突然
終	糹 冬
終於
船	舟 几 口
口	囗
答	⺮ 合
回答
禮	礻 豊
物	牛 勿
禮物
頭	豆 頁
頭發
關心
腳	月 卻
生氣
哭	吅 犬
畫	聿 田 一
輕	車 巠
年輕
包	勹 巳
腿	月 退
忘	亡 心
忘記
搬	扌 般
樓	木 婁
遇	辶 禺
遇到
聞	門 耳
新聞
較	車 交
比較
雙	雔 又
見面
經常
城	土 成
市	亠 巾
城市
一會兒
附	阝 付
附近
借	亻 昔
響	鄉 音
影響
認真
差	羊 工
銀	金 艮
行	彳 亍
銀行
安	宀 女
靜	青 爭
安靜
多麼
餓	飠 我
根	木 艮
據	扌 豦
根據
乎	㇒ 𠂇 丷
幾乎
後來
動物
一邊
舒	舍 予
舒服
般	舟 殳
一般
叔	尗 又
叔叔
疼	疒 冬
遲	辶 犀
遲到
歷	厤 止
史	中 乂
歷史
啤	口 卑
酒	氵 酉
啤酒
短	矢 豆
經過
周	田 口
末	木 一
周末
慣	忄 貫
習慣
園	囗 袁
公園
乾	龺 乞
淨	氵 爭
乾淨
鳥	白 ㇉ 一 灬
健	亻 建
康	广 隶
健康
樹	木 尌
糕	米 羔
蛋糕
元	二 儿
客人
議	言 義
會議
奶奶
褲	衤 庫
褲子
鄰	粦 阝
居	尸 古
鄰居
理	王 里
經理
層	尸 曾
燈	火 登
練	糹 柬
練習
爺	父 耶
爺爺
藍	艹 監
難過
中間
帽	巾 冒
帽子
司機
舊	艹 隹 臼
滿	氵 廿 巾 从 
滿意
騎	馬 奇
陽	阝 昜
太陽
極	木 亟
主	王 丶
主要
同事
鼻	自 畀
鼻子
角	⺈ 用
變	䜌 ⺙
化	亻 匕
變化
級	糹 及
年級
環	王 睘
境	土 竟
環境
胖	月 半
圖	囗 啚
地圖
面包
郵	垂 阝
電子郵件
耳	㔿 二
朵	几 木
耳朵
裙	衤 君
裙子
鮮	魚 羊
新鮮
放心
聊	耳 卯
聊天
南	十 冂 丷 干
熱情
卡	上 卜
信用卡
梯	木 弟
電梯
方便
洗手間
澡	氵 喿
洗澡
飲	飠 欠
料	米 斗
飲料
校長
平	干 丷
水平
業	丷 一 木
作業
襯	衤 親
衫	衤 彡
襯衫
績	糹 責
成績
碗	石 宛
阿	阝 可
姨	女 夷
阿姨
圖書館
文	亠 乂
文化
綠	糹 彔
掃	扌 帚
打掃
草	艹 早
冰	冫 水
箱	⺮ 相
冰箱
數	婁 ⺙
數學
自行車
急	刍 心
著急
瘦	疒 叟
提	扌 是
提高
起飛
矮	矢 委
鐵	金 土 戈 口 王
地鐵
育	亠 厶 月
體育
刻	亥 刂
護	言 蒦
護照
節日
盤	般 皿
盤子
一共
瓶	并 瓦
瓶子
街	行 圭
街道
鍛	金 段
煉	火 柬
鍛煉
感	咸 心
冒	冃 目
感冒
愛好
超	走 召
超市
月亮
飽	飠 包
有名
香	禾 日
蕉	艹 焦
香蕉
筆記本
夏	一  丶 目 夂
菜單
北方
網	糹 罔
上網
季	禾 子
季節
渴	氵 曷
燒	火 堯
發燒
不但
空	穴 工
調	言 周
空調
照相機
春	𡗗 日
傘	人 十 𠈌
斤	⺁ 丅
公斤
個子
熊	能 灬
熊貓
刷	尸 巾 刂
牙	一 ㇜ 亅 丿
刷牙
復	彳 复
復習
冬	夂 ⺀
假	亻 叚
請假
中文
秋	禾 火
句	勹 口
句子
李	木 子
行李箱
筷	⺮ 快
筷子
皮	丿 ㇆ 丨 ㇇ ㇏
鞋	革 圭
皮鞋
爬	爪 巴
山	丨 凵
爬山
板	木 反
黑板
趣	走 取
感興趣
詞	言 司
典	曲 八
詞典
留	卯 田
留學
颳	風 舌
風	几 䖝
颳風
黃	廿 一 田 八
河	氵 可
黃河
死	歹 匕
干	一 十
所有
許	言 午
也許
不過
發生
切	七 刀
一切
抱	扌 包
歉	兼 欠
抱歉
感覺
肯	止 月
肯定
棒	木 奉
以為
掉	扌 卓
活	氵 舌
生活
之	丶 ㇇ ㇝
任	亻 壬
何	亻 可
任何
與	臼 己 丨 一 八
弄	王 艹
卻	谷 卩
繼	糹 㡭
續	糹 賣
繼續
夠	多 句
父	八 乂
親	亲 見
父親
全	人 王
完全
可是
談	言 炎
好像
警	敬 言
察	宀 祭
警察
呀	口 牙
況	氵 兄
情況
只要
份	亻 分
底	广 氐
到底
成為
永	水 丶
永遠
安全
計	言 十
劃	畫 刂
計劃
倆	亻 兩
停	亻 亭
感謝
敢	一 丨 耳 ⺙
從來
贏	匸 丶 口 月 几 貝
消	氵 肖
消息
拉	扌 立
原	厂 白 小
原因
連	辶 車
確	石 隺
確實
挺	扌 廷
保	亻 呆
証	言 正
保証
受	爫 冖 又
接受
改	己 ⺙
改變
麻	广 林
煩	火 頁
麻煩
出現
管	⺮ 官
不管
甚	甘 匹
至	𠫓 土
甚至
保護
真正
結果
當時
至少
律	彳 聿
律師
演	氵 寅
表演
無	𠂉 卌 一 灬
猜	犭 青
咱	口 自
咱們
進行
內	入 冂
否	不 口
是否
調查
功	工 力
成功
慮	虍 思
考慮
約	糹 勺
約會
通	辶 甬
通過
開心
母	㇗ ㇆ ⺀ 一
母親
主意
倒	亻 到
釋	釆 睪
解釋
聯	耳 幺 丱
聯系
証明
命	亼 叩
生命
難道
由	二 丨 凵
指	扌 旨
危	⺈ 厄
險	阝 僉
危險
討	言 寸
厭	厂 猒
討厭
醒	酉 星
樣子
有趣
部	咅 阝
部分
理解
任務
使	亻 吏
轉	車 專
博	十 尃
士	十 一
博士
緊	臤 糸
緊張
棄	亠 厶 山 一 木
放棄
概	木 既
大概
重新
其中
來自
本來
並	䒑 业
並且
直接
對於
正常
遍	辶 扁
冷靜
方法
扔	扌 乃
能力
另	口 力
另外
鬆	髟 松
放鬆
丟	王 厶
負	⺈ 貝
責	龶 貝
負責
夢	艹 罒 冖 夕
戴	𢦏 異
誤	言 吴
錯誤
隨	阝 遀
隨便
經歷
支	十 又
持	扌 寺
支持
建	廴 聿
建議
則	貝 刂
否則
光	⺌ 兀
排	扌 非
安排
鑰	金 龠
匙	是 匕
鑰匙
信息
全部
首	䒑 自
首先
交	六 乂
台	厶 口
堅	臤 土
堅持
生意
即	白 匕 卩
即使
處	虍 処
到處
挂	扌 圭
道歉
憐	忄 粦
可憐
實在
騙	馬 扁
諒	言 京
原諒
亂	爫 龴 冂 厶 又 乚
差不多
研	石 开
究	穴 九
研究
擾	扌 憂
打擾
正確
收	丩 ⺙
秒	禾 少
同時
供	亻 共
提供
輸	車 俞
碼	石 馬
號碼
座	广 坐
比如
嚴	吅 厂 一 丨 耳 ⺙
嚴重
脫	月 兌
陪	阝 咅
法律
值	亻 直
值得
使用
方面
原來
論	言 侖
討論
說明
仍	亻 乃
仍然
動作
受到
趕	走 旱
懷	忄 褱
疑	匕 矢 龴 疋
懷疑
拒	扌 巨
絕	糹刀 巴
拒絕
演員
破	石 皮
此	止 匕
因此
案	安 木
答案
活動
既	白 匕 旡
既然
通知
不得不
無論
刀	㇆ 丿
適	辶 啇
合	亼 口
適合
失	夫 ㇒
失望
允	厶 儿
允許
意見
獲	犭 蒦
獲得
要是
邀	辶 敫
邀請
儘	亻 盡
儘管
浪	氵 良
費	弗 貝
浪費
敗	貝 ⺙
失敗
責任
美	羊 大
麗	丽 鹿
美麗
壓	厭 土
壓力
味	口 未
味道
厲	厂 萬
厲害
出發
奮	大 隹 田
興奮
觀	雚 見
眾	罒 亻 从
觀眾
反	⺁ 又
反對
精	米 青
彩	采 彡
精彩
感情
演出
愉	忄 俞
愉快
開玩笑
雜	亠 从 木 隹
志	士 心
雜志
合適
廣	广 黄
廣告
自然
深	氵 罙
取	耳 又
短信
地球
帥	𠂤 巾
推	扌 隹
鍵	金 建
關鍵
竟	音 儿
究竟
恐	巩 心
恐怕
躺	身 尚
聚	取 乑
聚會
方向
幸	土 丷 干
福	礻 畐
幸福
接著
技	扌 支
術	行 术
技術
困	囗 木
困難
正好
提醒
旅行
激	氵 敫
激動
驕	馬 喬
傲	亻 敖
驕傲
毛	㇒ 二 乚
許多
順	川 頁
利	禾 刂
順利
職	耳 音 戈
職業
賺	貝 兼
址	土 止
地址
於是
拾	扌 合
收拾
圍	囗 韋
周圍
愛情
尊	酋 寸
尊重
十分
授	扌 受
教授
超過
寄	宀 奇
順便
無聊
目的
低	亻 氐
剩	乘 刂
複	衤 复
複雜
社	礻 土
社會
故意
好處
竟然
示	二 小
表示
印	㇒ ㇗ 一 卩
象	⺈ 口 丨 豕
印象
出生
估	亻 古
估計
地點
輕鬆
作用
舉	臼 己 丨 一 八 二
伙	亻 火
小伙子
著名
免	⺈ 口 丨 乚
免費
傷	亻 丿 一 日 勹 ㇒
傷心
記者
仔	亻 子
細	糹 田
仔細
巧	工 丂
克	古 儿
巧克力
辣	辛 束
互	一 彑
互相
廁	广 則
廁所
程	禾 呈
過程
申	日 丨
申請
引	弓 丨
引起
展	 尸 龷 𠄌 丿 乀
發展
畢	田 一 二 丨 艹
畢業
式	弋 工
正式
廚	广 尌
廚房
專	十 日 丨 寸
專業
吸	口 及
吸引
心情
祝	礻 兄
賀	加 貝
祝賀
條件
千萬
糖	米 唐
趟	走 尚
由於
密	宀 心 丿 山
密碼
倍	亻 咅
擦	扌 察
尤	尢 丶
尤其
驗	馬 僉
經驗
盒	合 皿
盒子
乾杯
看法
髒	冂 ㇆ 月 艹 歹 匕 廾
藝	艹 土 八  丿 ㇈ 丶 二 厶
藝術
速	辶 束
度	广 廿 又
速度
勇	龴 男
勇敢
數字
暫	斬 日
暫時
優	亻 憂
秀	禾 乃
優秀
笑話
惜	忄 昔
可惜
省	少 目
笨	⺮ 本
科	禾 斗
科學
餐	歺 又 食
廳	广 聽
餐廳
各	夂 口
距	⻊ 巨
距離
窗	穴 囱
戶	丿 尸
窗戶
空氣
護士
悔	忄 每
後悔
大約
內容
規	夫 見
規定
效	交 ⺙
效果
金	全 丷
現金
童	立 里
兒童
篇	⺮ 扁
漫	氵 曼
浪漫
態	能 心
態度
自信
驚	敬 馬
吃驚
熟	孰 灬
悉	釆 心
熟悉
按	扌 安
按照
紀	糹 己
世紀
憶	忄 意
回憶
相同
重點
教育
受不了
膚	虍 胃
皮膚
區	匚 品
區別
左右
陽光
頁	丆 貝
章	立 早
文章
言	亠 二 口
語言
標	木 票
標準
管理
誤會
橋	木 喬
舉行
肚	月 土
肚子
僅	亻 堇
不僅
餅	飠 并
餅乾
際	阝 祭
國際
信心
抬	扌 台
競	竞
爭	爫 ⺕ 亅
競爭
湯	氵 昜
作家
誠	言 成
誠實
顧客
存	𠂇 仔
扮	扌 分
打扮
流	氵 㐬
交流
齡	齒 令
年齡
小說
符	⺮ 付
符合
交通
共同
稍	禾 肖
微	彳 山 ⺙ 一 几
稍微
增	土 曾
增加
敲	高 攴
適應
苦	艹 古
辛	立 十
辛苦
然而
耐	而 寸
耐心
將	爿 月 寸
將來
沙	氵 少
沙發
